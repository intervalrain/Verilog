`timescale 1ps/1ps
`include "lab1.v"

module moduleName (
    ports
);
    
endmodule