`timescale 1ps/1ps
`include "lab1.v"

module lab1_tb;

    reg x0;
    reg x1;
    reg x2;
    reg x3;
    reg x4;
    wire F;

    lab1 uut(
        .x0(x0),
        .x1(x1),
        .x2(x2),
        .x3(x3),
        .x4(x4),
        .F(F)
    );

    initial begin

    $dumpfile("lab1_tb.vcd");
    $dumpvars(0, lab1_tb);


    x0 = 0; x1 = 0; x2 = 0; x3 = 0; x4 = 0;
    #10;

    x0 = 0; x1 = 0; x2 = 0; x3 = 0; x4 = 1;
    #10;

    x0 = 0; x1 = 0; x2 = 0; x3 = 1; x4 = 0;
    #10;

    x0 = 0; x1 = 0; x2 = 0; x3 = 1; x4 = 1;
    #10;

    x0 = 0; x1 = 0; x2 = 1; x3 = 0; x4 = 0;
    #10;

    x0 = 0; x1 = 0; x2 = 1; x3 = 0; x4 = 1;
    #10;

    x0 = 0; x1 = 0; x2 = 1; x3 = 1; x4 = 0;
    #10;

    x0 = 0; x1 = 0; x2 = 1; x3 = 1; x4 = 1;
    #10;

    x0 = 0; x1 = 1; x2 = 0; x3 = 0; x4 = 0;
    #10;

    x0 = 0; x1 = 1; x2 = 0; x3 = 0; x4 = 1;
    #10;

    x0 = 0; x1 = 1; x2 = 0; x3 = 1; x4 = 0;
    #10;

    x0 = 0; x1 = 1; x2 = 0; x3 = 1; x4 = 1;
    #10;

    x0 = 0; x1 = 1; x2 = 1; x3 = 0; x4 = 0;
    #10;

    x0 = 0; x1 = 1; x2 = 1; x3 = 0; x4 = 1;
    #10;

    x0 = 0; x1 = 1; x2 = 1; x3 = 1; x4 = 0;
    #10;

    x0 = 0; x1 = 1; x2 = 1; x3 = 1; x4 = 1;
    #10;

    x0 = 1; x1 = 0; x2 = 0; x3 = 0; x4 = 0;
    #10;

    x0 = 1; x1 = 0; x2 = 0; x3 = 0; x4 = 1;
    #10;

    x0 = 1; x1 = 0; x2 = 0; x3 = 1; x4 = 0;
    #10;

    x0 = 1; x1 = 0; x2 = 0; x3 = 1; x4 = 1;
    #10;

    x0 = 1; x1 = 0; x2 = 1; x3 = 0; x4 = 0;
    #10;

    x0 = 1; x1 = 0; x2 = 1; x3 = 0; x4 = 1;
    #10;

    x0 = 1; x1 = 0; x2 = 1; x3 = 1; x4 = 0;
    #10;

    x0 = 1; x1 = 0; x2 = 1; x3 = 1; x4 = 1;
    #10;

    x0 = 1; x1 = 1; x2 = 0; x3 = 0; x4 = 0;
    #10;

    x0 = 1; x1 = 1; x2 = 0; x3 = 0; x4 = 1;
    #10;

    x0 = 1; x1 = 1; x2 = 0; x3 = 1; x4 = 0;
    #10;

    x0 = 1; x1 = 1; x2 = 0; x3 = 1; x4 = 1;
    #10;

    x0 = 1; x1 = 1; x2 = 1; x3 = 0; x4 = 0;
    #10;

    x0 = 1; x1 = 1; x2 = 1; x3 = 0; x4 = 1;
    #10;

    x0 = 1; x1 = 1; x2 = 1; x3 = 1; x4 = 0;
    #10;

    x0 = 1; x1 = 1; x2 = 1; x3 = 1; x4 = 1;
    #10;

    $display("Test complete");
end

endmodule